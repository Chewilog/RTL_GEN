entity SignedTest1 is
    port(in1: in unsigned(3 downto 0);
    out1 : out unsigned(3 downto 0));
end SignedTest1;